�`  =��N����9+fo�x�       c ��x ' }���.   � A�    �> ,  �   
�#<� 	  �� 2 2  �   � �{ |� { . z lv { t }z�}'� |�{ }�u|',z y uz't lm z��
ll t	�l�| tdtl tl�d�t���| 2 tdl
�t�t uy�l�dtt*$���d�||%l��|�
dl
��� �t	ey�1��|	�|d	(�tt1l�d|�tl| |l�	l||ld,< ���,� t|t��C��tl ||( �tl| l l� �Pt�� �ld�ttt*Lll �| |�t l/,(l�d,� v,{ �6t( t	�l�l	�*� ||�dm|�l�Tdl�ddl
��|�d|l *D lll|�t �|t	tl l( �|l( t%|t,����t t}%}�|d| �ldddl l||
| d�"l�pddtt| �l|t��fy t
�l�l|dll
|(t (� |l| �� |� �tl|| �	|!d�tltd� ��l�d��� tt� ��|�d|&� �t �
t |	�t��ltl�td(D |�ld(ltt��
��d(� l� *� d*��ltdd�t �,�tl�t�t d� �d	�����l*< d�d� lt|!�� �t �Zd�� (< �|�d�t l �d�||, ttl| t| l lt| �*� tl �|td| (� �t l l�$dttv��� l�� |ll l�l� dllldlt| �ddl �|tl l( lt�lt|3l|ld| |�
|!�d� (� d|(||dtdll| l l||(� d(|� |�|tl �d* l��lt
���	lt| �t�dd�d�����t�� dl �( t� �(��tl�d|�t�(� d� t �� �lll�lll�|#���|�(\�|��|,$ �� �� l�ddd||l ||tj��$t�|l lldll	llll� d�|�� |���l4tddldl
l�t��l�l0l td*l�dll�dl ���d* |(< tl || ��l�d|�0ddl0d t|�"�!l|� ,�d��
(� �td
l l|l�t�|�� t(, |dtl ���tt� l
dOld�-,$|7t	l ����d
t	(� �lt���G�t lll* l� ��	�l��d* tl(d"D!�|d��� �( t*d |l"���dtl�* td| || l l� �l|| �l
$D(��(�td|t| t"�9(d7tt| � �t || ,| *�dld�� tl� d.l|*4�dt�� �t l� �
�ld|� dtl dtd�Ktd�tlD��� (L �| � (|�t dd� d�dtl tdBl�� d�l�����
*\ td�|ll|�|�lllll t�tt&��d(� �0t|�
dl �t |� dd
l	t
�d�
d"<9| *t |�dd��d�dl �&d|�| ||��|�|�|� (|�(� ��t�dll	tl�l(Tt�� l�|d(� |	dl t�tl (� |�*L ��l|�t(4l�d
tll �	|l� td�llt* l�|"||��� (T d�lddl t�dl �|�dt��d��dt|�dl �* ���l�|�|�| dl� | (�|g�t
��|'ll ll |��2�l|��| ��l
�� �	l�dt| l �tl�tl dd	|
�tl d�t * dl �d� tdll
||l(\ dddl d|t��Bt�	ll |��|d(� |'�l�t�|� td| dt(�t(T|d|t��d�dld
l( �lt��Hl	�I�l*��lll l���tl
||l �� (D �t (� |(D (� lt�d� �l�|"�,�tl (4 t
� tlt�|( d�1��$lt
| � ��|l �Dd��dl |�z�||&(l �
dl �|$�&dt�|�t�| |l(| dt"�Q���|�dl d| l	l d| dC� ll �l|,� tU�dt(4 �	|� t dl �� l�t ��� (� d�l|ldll�t	|dt|dd|l�d
��	d�� |dll�|t|	t.� l�dl ���(< *�tl
t| l |	|l�lt(T �t||��U|�t�l"dt� |d�(� t�l*� ��|Dd��d4l |(� �l	t|l!t|l||l| , t(� �||�(�
��� tt| �d� |	t||�td	d* tl	d�l��d|	�l|� tdl ld�| ( �dl�t4L(� dtdt*, �(� dt
dt( �Il�t�-l|| ����l|�tl	��t �� ��t� |dl |N���dtld�t�d5d�dd(� ��dtlll� d|| l dl ��,| ���t�(< t	� f} �t|l_�tdl td$*l��lt�Mdl"d<��l�* *, �t t* (��l>lt"d�� |�ll
�* t, ll t���d� d�"�"�|l� ,��lplt| l �lI|�	��tl dd� �t � td0���� ddtd|l d|�ll �|l |dd� tllt
|d�ldk|l|( td���|tl ddd||l(Ldl �dl �d�d�|�tl tl
| ldl ��(� dtd��8�_tl	ld| |d���t�l����tdtw| l ��|�|dd�ld|| tl� d(���dt|| t
|� ll�|�, �lt� * |	�l��| ll �d�llll |
� |tl d|�5|�lt*ld� |Xd|� |l ��| �	�	t�ll �d�d�d�"�E(���l� ����U�( t�d	t(� �� (� l�| l ��dtd�d(($ tl �t8d|��t|| dltll l|� tl �t��d!||� |||dl |d� tt| d|d|� ddl
d| �dt|
� �| t�|� �t
d����|l� �d
l �|dl �dVdltd||| "�7tt	| ll|| l (L d|t| � �tl| � �t	|| dt| ���t�|||tl	�tll��d
��|dtltl �tttl �t �t $�Dt�ldl �t lI��
ldl |l� t�td��tl�~�ltl l�t d�t� *< |	t| �t �@��| d| |/tl( ddl�|d| �d|| dtl�d�rd|	l �l� �Rd��|�� l�%���� �l�ddl �� d�*� ll �|��dt4 ll |(� �d�(� lt�d� (� l�����t(� �ld� ��|� �l�|'.��d�d� �l�lldll t|l ll�, ddtl tl l�d�lttlll|�ltl�t t�Rt dr�� ��tt� dl |dd� tl �l�| �t� |d
�dtl� |(T �l��	�(< d��l��(L�td| l �tl
l ll* t�ll dl�ll dlt�d|| � |l	(T dld<dlt	t��
lt��t�td|d�t��tld(��|�| |�ll|�|l || � |�t l"�5��|t��t��lt| d.|l�d�l	�|� dl ���� �l�Ӵ��ttt��	t |t�g���	tt��d|lt�t (�t(� d� l	|| �tl �|�lt�|lllltl| |l ||tl��|� ��� �|l	��	(l �ll�t||ll �dl �*T d|��t���|l� tl �d�&t�lll t|� |tdt|l l�dd�tdtl �dtt(t ltl ��, �d|ll
(d�|�� �d�l|�tdl �|*\dl �#|t���� lt
|l |l||��|�tt| � �| |tl|l���dl t� td| l|l� �|tdl t� tl�d�lttl"d�l� ,�d�dll�t tl �dtdl* ���ll��t l�Kd�t tdl|| "�*l�
| � �l�||| � |l �l
l |(\��	|ll!��l�t(4 ���d
�d��dl ��t-�| t|ll d| l t	l *� ��l|| � l�tl l|l| |t@�|��(, �|d�l��	|�|'dl *, ||�%tl tll��t
|� ����l
|��dl� �t|d| t�tdl tl l� 0 ||� (*� |�| |lt	t&ll| l �t l d� *< �'ld
d���lll|llt�$Ndt��dd�t|l� �|	dt|�d��ll4t� dl�|�|l�t� �t�l�(T l|l t�tt�tt.� �t|t|| �| |l�d�ll dl ��tl (d ($ �dl t� |l *T�dt/tltt��| �l�� t�l	�lll|9(�>dlt.ll |( dd| �'l	d| �%�ttt� |�tl"��ll l| �ld0 ltd�f�d�dl �dddl|t( *D (�|||l| l �d
t(� dl�	ld�tl d�|�l��|td|l��� dd���tt#"�r",Etl |�dt� �	l�� |�d|��lddt
ll�� |�� |� t �O�|d(� ���t� �m}%ğd|Zll �	( dt| dl�>tl �dl| l ll t|| �"dtt�|l�d�|�l$<$����l
ltt	tl| �| t	|l dl�*4��dt�. |t*� �<�|t� d|���|�t �d|�t�|t��t ���&�dt8dtlld(� �"d=d��(� |� �| t| �d ��|:�
|�|��|(|l	(� t�(<�td.� d�dt| �t^*� t��t ���l/|ddl$t,�|�ll l| (� t(� |||(l�� �|� �l�d�����l|�, �l�|	��||�|l l|�(d(l dddt
� t �|d� �l|�	ll tl �dl| l| |��
ll l�|��(� ll�ldl (, dl t|� t d| *�(� ����� (�� l�t ( |�l	d�dl �lt||plt| �t d�	�lt�d|| �	�lll lll�Ť|(d��Kd��td���dl�td| l |�t d|�l� �,� ��|��|� "�%l
ddll ��|��d�|	l�ll dl || d� t (T t��!d�"�Xl����|�ll ���� ���'t
�|tl l|l�| |� l�ltdlt|(t|d	� �ld�l�ltl l��t |�ddd����t �
�dQd�( ldl� d|d� d�-dll |�tl �t l��� l
l| tt|( l�l|�dt|�l,l |d|t���d�dt� tt	| � t�/�� |	d|l�� t�
|,t�d,� �dl �($ ��	�� �xt
d�d|| �dl(�dl �|�� t,t |
�l4�( �t (� ll���d�*|t�dl dl� �*�(Tl�d�(< t�	t �	�'ll��Ctdll l� |l|"�(ld� t �t l*�$&tdl |��(T �ldt|| (L t�t� 	$ �`t�|�(�
� tdttt�td��|ȴt ��t , �ll2|	dtt	|�tl dtt�d��tl��	�|l ,< t|lt� ��	�d|�d,��d"(�*T l|l �d
|( lt�td� dlt��l�t t%l ��|� ��td
,$�l(d t(� l|!l l� dkd.\ d�	��ll���tdt�|*� |	|l |ll|l|l ||| �|d| l(��||tl |l&ll �t	d�?��tdl l| l d	| l� � t��l� lddt(T �l� ($�l�t �� ttd(, d�l�l($dd|d	ll�t�|ll |l �ll �t �|l	ld|l�dtt�tl� dld�;|ll�t l��l�|d|�l||� dt�� (L �d�|�d	l t�&<C|t| l| �d� ��d#�| �t ,|l�| tl (ll|l || dl d|� l|t
�d�d�|�t �*L �t&tt�td�t l �d���t�<d|� t |�d	(L ��|t��t d�l*� (\ dt!dt| �t �d�|t� |(�d�	dl��ll |d(|��l)dd� |l �tdt| ���t ��t	ll |l ��dl &�%d|dl |d,|4�t���,� *�|l#d
�t tl �	�d"�||l d�d �|ttl ltl�t $�?�
�ddl dd	ll d|l *ldll|�l|�d�
|l|l|l �| |� tl ddl |tl� �� l(d |�| t���l
|l� �	|�(���|��(� ttd	||(� |�"�+ddt�(� |l	tl �tlltdl d	|| ll dp�ll(,�ll|l�I��t ||l
|l| l�� (��(� ��� dt�	� |��|t�0�t�tt, ||| � �� l�
l|� ����( |ltl
| |l l|�dl �d
lttl(\l	ddt�|* �(D |4� l�|$�K($�;",Kt�(� �|d|*�|�l|�|l t	l|| �*, |l �dd ( |�|	��W�ll| �� �d|l ��
|
lt#l�t d���d�(� d�d|( |�d(� t|t"d� l'l|�� t� (D ld|�� t��l�ddl� t��l���t|�l|��llt
�d� td� l
|� � t� (D "4�t
d| ll�� l
�2�tt�t|�(L �dl �t	|tdt�t|
�t �N"l*ld�t�dldl || l� �� �l���l��l"#�ddl*���t l �d( �tl ��||�� ����tt�|l�l�t&dl ��(� l�l��t||	��ttd��� l(� |k�,t�9|	ldld	� ���,\��d
l4tl
dt�t�d
t|dl� � |l| || d��tdt.� ||| �t� |dld	t�tldt|dl l�l0L d��||l� d�tldlt� dl td(, dd, �l����� t�ll�d� |�8ll��| ltl| �t*|t�&�>�2� t|ll d� �!(��Jtd
�d� �d��l|��dl�dl t� ldC� t �7�( �dll�*�@�l|t5�|
� ll��� tl d�dd�ll�%|, td��|ltlt�(4 d|(D t,4 l||�l,<���dt� tt| ��(t |l	d| || t� dt�t�
l �|� (� �d	( �ddtl| l�	dtt|ll*� t|ll �d� d	l dD|� �| |�� t ll| |l l|l (� d(4 lt�l�d|||||�d��dll t|||l || �l���( �|(tl tl l��t����tt|�t� d�|d| �d�d� dl ll t(t�|����dl d| |l� �(� ��� &�&t��lllt(\�|l ��9�tt� .�||
���| |tl�(tdl tt� �|�
��l	|� |l (4 ���. dl �&*tt�*�d��|	($ t"�&ttdl �	d|����d�
t � l|���"\"l|�t �dl |����l�|� *|�� dt|l ||, �� (4�t�(D�ddl|��l(,dt.D �� �d|||l ll�t tl �� t,tdd�|��(, l$A�(� |(�|d�(�|�|$� t|�d* tl �t �t |tl lll|�dl ||ld��t ��ld|��ldl� t |tt� |,� �l�|t| ttl �d( �e���dd't||dt�td	td(�lddt| ��l�ditd|tll �tl tt| �ll.� ||�d(�(l |(� |tt��t,t |l |�t d�t l dl t|�|	tt(, d��*�/|itd�tdt-l��| (� d���ddt'| |d�|�t d
tt�dFt�lll d|l� tdt�td� l��tll t�dd�t�� |t2d,� �t �d���( |� |
*���	td| *�l|ll l�
���;ltl ��dll �( tt����td/� * l� ���(4 d�dd����l�t�d|dl ��(� l||�l��t%l�d�d�	dl �|l ���| l ��d��dlt�t �B|Mll, td| "�Q�td��|	�|dl l�
|d| tll!�| (�l(D lt�|l|* l���lld(��|ll	�l�tl���|�d|� |*|l��|t(��|�dt|tllll| ��tdldd��	ld	|��|l| lt��|	d�tddt�t�|d| t�ld(� dd. |�
dld*d	t||d� l||��t t	l�dt� td
t"L8| *� |�| �||
d��d� �|t	tl l(| �l�ldd�	d� �	��| �#d� ��dd(� |�l� �(� �� �"��(� �	dl |d||l� |d�	�tl
�� �d� * l( ��t	lt�ddl ll lt	� ddd"/t�|"l|l�dd� t(� l�| "�5t�* l
�l|�d
d|� |
d� ��*��|dlCdtl|�dl �	| � � | l| d|(< �t���d�tl�t�*d���lt��|d� ���
ll dl l(\|	�( dltl�* |tll (� tl dtl�|�|t(< d��|�|dl |�(4	���| (Ltt(D |�|� |��tl��l* d|��ld� t
l t| tQ�|ddt| l| �����0 �|� �9||� t�|l ll (� l�	|ll dd�t�ll
,d tl ��t(t|* d�� l�� t"<5�t(�ll d|l|��|l �)dl �t t|l. *�|d
���||t�*$ dtdd*l�=�|� ��lC(���"�=|�|t�	d( �l|�ldd�d�dtd0L d(� �l�d�tt"�Pdl lt� t d�� ��t
l�"�<�t�	d�d	t�lt(< d�'t�dl�l( (L �Ml1l�(�t|dl���l�|l ���|�t ll *, lt��|l( �
|�d��t t| l �t��d|t
l ll �t� tdtlt(L |	�d�|tl� ���, dl (T �	*< d�|���l�||�|d�dt��|Zt( d(4 �d|d
ll ��t |�tdd�|� �|`l�t#t���Ztl�t |	tlt� �t l���l|d., llll|�ll |�dl�t� tl��lt(� �|�� * tl l||d( tt� l( l|�t*<�l�dll |	�d�
|ld�t�ldd�
d�lK|����d
�dl(�dl��t || �d�t� ltt	| l ll d�tl �|t� t|||., l(� (� |dt
| |� �ld|l |( �� � �ll t�d	($ l�� ,D l!�d|�|t
�ll0� �|dt�d�|ddll|�t l d|7�� t
�|�l� ����� tll� dll d| �|�dl| �dl tl�|*� ||�|9�t|� |l tl| �(�d�|'tftl|
&�$|� |�t�� �d(�t d	t
l (D*d lt|t1� ll��t|t���ld(L|�� dl| d ����t l tll|�td���dl��ddl�t� ��ttl �|��� d	�d(| l�* |d	|���� |�l� t. d>dtl
t	(� dt� � �(� ,< ��dl��d	dtl |�( lt| $Dtt� td�d(��t �	�ll	� lt
��|�,�| l;� �� t�t(	l�dt���|dll *,�t��tl t| ( t|	d| |l� ��ttl(lt� tl d��|�� �* �
� t�t l d( ll �l�d�d""4%d"�'��|
d	� dl tt,t "�Dlt�tl �� dl t�|*�|l �l��|l�i�|��|d(4 ll �ld
|ll ��|*\ ||t��tt�tl|| d| |t� td�|�� d
l|d�dl�l(Tltl l� �ll �| �d� |�+(�ddl�dt
llltK��t|tdd||�ll|d
l �ll |l�
lll �� ddd| * l�td�(� ��|l |l l(��l�ll� *$ tl �|��||d*\ ld|�� �� ���|Td�(� �t	l ����t|#|��lt� ll�dl t|�d�d	�|t|l l. tld
t|�d
l|l�� ll
t�tt
d�$'t�* dd|| l�tl �| l ll	l �t tt|�ll �	t� (D tl| t�tdtlt�|l l|l �,� |l||��|l�dt�d�d���t,< �t�l�ld�t� |l t�| � �l|* |3��tt�� �d�t lt��dl |� �(� |�tt���ll �
ll �(tlt� d��|� dH||l |d� dl
� l(� tl t� d
|� t |�	d	ld	� �,� t.llll|� d���	(4 t���|�� ��||t�d��t tl l�l�|l l�tl d�
�| �0(�,\���(<'��t�dl �d���||� ll |�;�� t��t�|��l�| ��|������ dlt�ll ��|�tl d| ���t���d|l �d��	� t��( l�td� * tl l|� *� tt( |(\t|dl ll�tt�$$�d2d||�d( �$<&�|�� dt(� �l�	�t�ddd$l4d�� (t �d�3�lld| tdd�t�|� �|t�ddt�stdl� �d��	(t d��t��tdt�| �ltd��t�t���t �tt�
t d| �l�|� ||���6dl �d|(4 d� d	��l,D .4 |� �d|ntdlt�|l�� ��tl |!|l ll*||Yl|l �ddl d�tT�d* lll";�tdtt� t ���tl� "���ddt| ��dltdl ��
dl �| t||l ��ll| �� |(� d|tdd�|. $D��|;��||��l�(l|d)l|d�ll |l �ll ��d	l*$*, �ltd�dl ��ldl�t� d���0 *| ��tl��Cl� d|�|����td��t�d/l	t�, ll |	l �l�ll� dl �|l?��ll ll� dsdd��� ldl |��
td( |t�d� l��t tl d���td�lt�|.|l lt�d� �
t�, �.\*� |
d��l�td*4 |d� lt(� ���-�ddt&$Q|�� l,\ �|*�d�|��t l""||�,� l|l (��l
,� tt�td�*|	|t|��t���|d��tl�(t �|���t l �ldl ��dt� l
l t|l lt}�	��t��t ��||
�(� �d� �tl tl (� t(�t�dt� t	|t�t�l|t%d+d�� �"ll �l�| |�	ttdd|dl |��� l|t�t dd� ||l�t	lddll l|| *� ll d���l|� d
�t |
l "L"ll��tl d��|�d(� dl ,��t l ll l|| l	� �
tl �d
dl, �}��dt�ll
*< ��	lddt||t
|lld	d�lll d�dttd
|������d	t��� d�d|�� ,� ��|
���lM|�l�ldll�|(� tdkt(T ld	�t(l l
tl( ddt�l�t * l||t	|| ��|�dd�	|�l�� d��l|$�|l	�l����� |(��t|� d(� "$&t�t|��"�+�d�||l l���d	|dl ll lt*| |l �d�t�(�ddl ���B��l� dd��|�d� �tl�t �ll|� �t|l ��|�ddt| (� �	d�t� (T ��� �%�� |l� �!ll (t ���t	ll (� ����( d�d�d�(S(� d*� tlt�t. |[dt�| t|d||l| � �|���Jlt
tt
|d| � �|d| |�� |� |� ���* t�|� �
|#�(|tdld6| �| �G�t�t�� ��td��dl �|�t l ddl��ll| ld|| |�|l lt�d
�tl��ld�d��|*�	|ddld|ll �tdd(�Y��dldd(, d�|l d�|��| �l. l||l| d�| l l�d�t ll l� ,4 ��(���
dW|�tl |/l!| tP��$�Ot(,�	ld�d�|(�tl|
t(< *� �*�(td't��l��0 �	d|���tl �ll�tt� t |�ldtdtll� 0 d�l ttlZ|dt|dU| ��dl d�t���"A���.�t�t	�l�|l t| l �d�| tt�l	�t �l|t�t�tldt| d| 0l l(� �lt	���Tt�,��	��ll �
�( dl�dctdl �tt�|tl�(�(� �t�l�(� |�d
t�I�(� tt� |ld$>|d�(d|d
l |�t �d. �tl�l�ldlll t�tdt�l� |l |�ldl ttdtt|| l� �� ��t�l�d|dt��d�l�|��^dl t| l �� (< *��	��|d"��l6td|| �
|�tl	dl�lt
��|	�* �ll*<l|t��(d ��|l�t ||l dl�|l (< �ldl�|�t ��|ld� |�l|� t |� t|l l��� �t|�d�t ll� l*�|d�ll t�t|�
t ll|� t l �l� l�d�
l�dl|*t���ld�*� �|�dl �|��d�t dl �. dl(� td* tt	(L tc|dl �*, �d�|( �|l�t �t�t ��tl7ll� ll d l| �t|| �tl�
t�d�(� d�tldl �t �l*| �|�
ll||�| �"4A|	l t| l� �d�	�tl l�Mt� �
|tl l| l �|t||l||�t�	||l t|� ����t �� ,�$�� t�d�l
($ tltl��t�l($ (� |l( �d�| � |( ���t�ttt�| tll	�-tl t|�(, �t!l�	t�lt� �	(t |l| tdl�t t| *|�l
d| (� �(\ �|� 2ld��l�| tl ��tl ld,T ��,d d
��ltlll	d(� �� ddl l"�� dl l( ��3�tl l| t�dl l��dl |�tl l�lt( �
�d��� t|�ll �|��ll �t l d��td�tl t	tl (�t"�5�� �tl �
|� l	� �dl�$)���t d| t�*4 t�%|� ��t tl |"D7�t����t
d( ��tt t�(� �
� t. �� ��*� d*< dl	|� d�|t4|l �t t(� ���l||l |	dY|� ||lldl|( �l(L *$ d*� ��t |$"*�|tl �t t� |d� � t=ltll �d|
� t �t(� ll	d.| ��
�ll�|t�� tl| �(tlll ll|l	�t�ldd�%��.�t�d�
��l�dq�ttt��l�t�( �dt
l( ���l�l���|�d�*$ d�l(, tl t��ll |d�d	� (T �	|l|��� �	|�|�
"��dl |&�h||l� t ��d�ldl�(d |tl|||l� �l�ddt� �d� l�|dj|(D |(4 t�dFd�t
ld�dtl t�td
dltl t| l |,l �d�dt�ll |dtl |�t, tlt��tt| �|"�|tl,| t���l	ttl��� d|t�ddt�(� ($ �t|�d|���| ��td"�=tll �	��( ��ldtl �td�(�t�t�d�d|����� (D t�
(T �l�t�t|l ,\|(�� |�	|d| tl l�t (�*\ |�l|�|��|�tl l!d*| �tl|	l�| �|	td� ������
�dd'� �d($ |	dl ld� d( t� ltt|
|� l(D |�($ �� t ||lt
|���t$�#|tl dll���ldl �	*� tl �_(d t(�Q�|d�tl1lt| tol�ddt� l�(� |	�l�l|t|� �|�*, �(D �d*� �|$�0|t�l�(< (Tt�t�|lltl	l |, tl ��d�|�l( �t
��(($ ��� �lt| � �l
�� �t d� |�ll|d|lG�| t(,�|�t dl t����t�t l (\ l�ddld�|� ��d� ����=l�d�d��� (d � d��|�td�|l?.�|(ttdd��� t� �dd(ld�($ �|�t ll lt| l l�dl�)l�t ��� dt| |l l( �|ld� d�d�t ld||�t�t� ltl��d� tlll| |�l�| ||l l| |�t*� ���dt��
l|t� � (� dt| (� d(��t (� ����l�dt| �|d� �ddt�F��| lt|�d|t�|t|lt0 d�(� d|el��t�d|�8 ��ll �"�!,�|
��t �dltl| ��tl!d( ltl| l��l|l l"T6�����t |
l||ll|��l|�t �ld| (T d�|�� ��ttt|l��*, �8dl t�0 tl (d tl�|||l�(� l(L �dl l>l|�dl	dd(t���| t| d�$�at|$\cd�l�ll �| |�|dd	0 |t� l���(| dl| ���ld�� �t �!dl�$�t �t t��	( dl �t
�,� .\ l.� t�|�� (t�|
0� d�dtl ll �dt	��l|�l�*L ���|���dl td�t||l (� t�l��l���ddl d� d��tl dl �dldl| || |l� �� ||� �|dg"�#l�t �d|��t�	dl/|l| �| l
���l)�|�(� |l �� |l |
� ll||d
�lt-| ll �|	dtl d|dl||l �l||$45dl( d�l�	dll ��t ( �|�l��
tl ����� l�dt�t t
d��l��l� � |(l��(Ttt��t l�l�| t	||lll|lll l| ��� �|t.|l ��td���ll |( �dt��l!|ll�t�tdtl d� �� ��dt� l
d� �tl �l�*, d�d�t��ll�ltt� l�t l| l |t�t�tl dt�( dt| l l|d
llll( ttdt� ���F�dtt�|d||�|���� t l |�
"Ԟt	�t �
|ddd� �|*ld* ||l �!l(�t |||
| l|t*�|ll �t (� ld|�� (|d�tl tll| ld	|�tdd��d�(t d�l�dt(� t� ||l l
| ����	�� |t| ����| �(� d�� ��l� tt�|ldl |d�dl .�tt� "�+��$ �� t�d|*Lt�dl tl *��dl |�Jdl tl (Ddd� tlt|�1�*<�tdd|*\�( ��	(� �(D dl�"�!��	t�* t�	l���d�$�#(� �*�����tt|�| || l ||�t|l� td��, �l�d� �d�t � ll| l �(� ��d|| (� (���	��t�� d@l|
| l ltl. l�
,d |!||2� ��t�� lt�t �|�	d|t,\�dl ��
l8l �|�|��*L ��|�(\|t� ld�dl�t|l lll|t
t�t��$<Mt||�d� t ||l	ll �||�� |�d
l tlt� tmt�ddl �| |tL�d�d�|dt|t|� l���dlttl l� ddt� | t| d� d|� ldtt�|+l �t�|�l�� dl t�	d�t|	|� ||)d0d�dt�l��
�,\lld|�t l�ll�ddt|l|$9t�l�,L ����9ltl l�,4�|tl t� tut��dt��d
|(\ t� �ll�dd�(, ���ll �� t�dt(� dl ��|dtl�+ddl �lddWlt(l tl �d���tl �l%��h��|t
|l*t ll	| l l|�t ��� �%�l���t�
ddd`l dtl!� ddd�d�M�(l |� �t ,| t,T �|l |ttl l, �||t* ��l
� �t�d(T (l(4 d�l�� ||� t
�� �Jtl t� ddl lF�(Ddld
� � �.\ �d	d*�:*Tl�'�l|(l�l�t ||��ddt*D d�|d�(� �t tdll	d�ldl| �d��{��� tt
(< ttll	l t	���dd���l� d|	�|l�t ��|( *�dt�	lt� ddl�	� �ttt| t| (< d|llld� t��|l�l( t�|�(t �t��d�	�*� d|l�t*l �lld| (ttl tt| l �"%ld| �|l td
�l*\�d( �k$� �dtl �	� d d�|t� t�ltd� dld��� �| �
|t|
t|� �t�|�lt��l|#|� �tt�|d,�lltl d,� tttld� t� ���	d�dl|d�| �
� ttdl$t&�d�| t� dl t�l��dd
���t�� ,d �� �	d�d
($ ttt� �
� �(� tt	� �	|l�| tlt
|(ttt�t+|l	�llt� l*� d%d|(� �|lt| � ��t�5�tl| ( lt�l��|l� .�ldl t��t �|$�t �
|t|�t�$��"��t ���t�(� d|
l t||�t td||
��|�||td| ���ll d* d||	d"�(l|| |||d��d� � d�t�l|�l�|l	l�(D t��d�l� �ll �� ��tlll�ll��l� t tl ��ldl l|| �	�|*l�l|�dl tl �|l �d. |l
t:t�|ldl|| l|�( ll(D dd,dl ��
d	|( ��|��|(� �| *| tHd,���dQ�	t�� ll| dl� t � ��ll d,\|l ddh��|dl| �t��*�l��d�all |��t	t
||( dl�
td||l	�d��lt|d��|��*4 "�&l	�|tt� d
�ll |�t�&4`|lt�( ��l0l�d�|	l �l�dl �t ltdl�� d�tddMll ���l�	��l|��ll l(�dt��t �t�d*� �t t|(|l|l��|dd|t	|�9dtd| t| t��'ll�"�ttl t� l"�@�|�t�d	t� ll l*Lt(� �	t|,\t�|D��dttd
dl |�ddd���|��*| l�l|1tl|	�| l t	�ltllll�|l|�t*t �d
l�� (� ���( �� t�ll |��d�)�	�t �3|��l1��l�tll� �l
� ||| l| �dd� �t|�l||lt��| �td���t�9�
|dtd|�dd( "|#�ddl �t ttd|l |�tl ���!� d�dl �	t(4 t	t�dl�($ ���ldl l(,t���|}l|
|�l�tl lt�l
d�tl� |l �ld|�l|�&�#t|�t�|� l	d�|� |�l�t t*d|� dl|�l|�l�(� l|t� ��tl ����� � *� l�,� �t=|d(� d��dl� ���
��|��td|dtd|d| tl |�|l ��d	�lt| (� ,�l||�dl ll d�l[�|td�| ltl |��d��t��d�dl�l�d�d�	( d�
t� �
td|�ttl�t|t(T��l|l l�ddl |tl ||��d|t| |ll ���( �|d� ,| tl dl �� |l ll*�t�d��t�|d| �l�*Dtd
*ttl ll�tE(�||t|l �?||����t|tt�tll�|d�  z | z | | | { { { {   